// Copyright 2025 Tim Tremetsberger
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE−2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

/*
  Testbench für seg_driver (rein kombinational)
  - prüft Einzel-Segment-Aktivierung A..F, G bleibt 0
*/

`timescale 1ns/1ns

`include "seg_driver.v"  // sicherstellen, dass Dateiname so heißt

module seg_driver_tb;

  reg  [2:0] pos_i = 3'd0;
  wire [6:0] seg_o;

  seg_driver dut (
    .pos_i(pos_i),
    .seg_o(seg_o)
  );

  initial begin
    $dumpfile("seg_driver_tb.vcd");
    $dumpvars;

    /* verilator lint_off STMTDLY */
    // pos 0..5 → jeweils genau ein Segment (A..F)
    repeat (6) begin
      #50 pos_i = pos_i + 1;
    end

    // pos 6/7 → default 0
    #50 pos_i = 3'd6;
    #50 pos_i = 3'd7;

    $finish;
    /* verilator lint_on STMTDLY */
  end
endmodule
